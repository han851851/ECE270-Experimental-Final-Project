//top wrapper, connects pong module's signals to actual pins on the pico

module top(

)

endmodule